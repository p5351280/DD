  module first;

  initial
    begin
      $display("\n Hello Kitty!");
      $finish ;
    end

  endmodule